module Replicater_8B (a, z);
    input a;
    output[7:0] z;

    assign z[0] = a;
    assign z[1] = a;
    assign z[2] = a;
    assign z[3] = a;
    assign z[4] = a;
    assign z[5] = a;
    assign z[6] = a;
    assign z[7] = a;
    

endmodule